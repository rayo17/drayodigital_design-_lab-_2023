module ShiftBit (
		input logic In,
		output logic Out);
		
assign Out = In;
		
		
endmodule