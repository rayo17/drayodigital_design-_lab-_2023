// Copyright (C) 2022  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 22.1std.0 Build 915 10/25/2022 SC Lite Edition
// Created on Mon Oct  2 17:18:14 2023

// synthesis message_off 10175

`timescale 1ns/1ns

module tareaFSM (
    input clock, input reset, input M, input [7:0] contadorCLK, input [7:0] contadorMante,
    output [7:0] registro);

    enum int unsigned { S0=0, Mante=1, E=2 } fstate, reg_fstate;

    always_ff @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always_comb begin
        if (reset) begin
            reg_fstate <= S0;
            registro <= 8'b00000000;
        end
        else begin
            registro <= 8'b00000000;
            case (fstate)
                S0: begin
                    if (M)
                        reg_fstate <= Mante;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S0;

                    registro <= 8'b11111111;
                end
                Mante: begin
                    if (M)
                        reg_fstate <= Mante;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= Mante;

                    if (((contadorMante[7:0] == 8'b00000001) & (contadorCLK[7:0] == 8'b11001000)))
                        registro <= 8'b00000001;
                    else if (((contadorMante[7:0] == 8'b00000010) & (contadorCLK[7:0] == 8'b11001000)))
                        registro <= 8'b00000010;
                    else if (((contadorMante[7:0] == 8'b00000011) & (contadorCLK[7:0] == 8'b11001000)))
                        registro <= 8'b00000011;
                    else if (((contadorMante[7:0] == 8'b00000100) & (contadorCLK[7:0] == 8'b11001000)))
                        registro <= 8'b00000100;
                    else if (((contadorMante[7:0] == 8'b00000101) & (contadorCLK[7:0] == 8'b11001000)))
                        registro <= 8'b00000101;
                    else if (((contadorMante[7:0] == 8'b00000110) & (contadorCLK[7:0] == 8'b11001000)))
                        registro <= 8'b00000110;
                    else if (((contadorMante[7:0] == 8'b00000111) & (contadorCLK[7:0] == 8'b11001000)))
                        registro <= 8'b00000111;
                    else if (((contadorMante[7:0] == 8'b00001000) & (contadorCLK[7:0] == 8'b11001000)))
                        registro <= 8'b00001000;
                    else if (((contadorMante[7:0] == 8'b00001001) & (contadorCLK[7:0] == 8'b11001000)))
                        registro <= 8'b00001001;
                    // Inserting 'else' block to prevent latch inference
                    else
                        registro <= 8'b00000000;
                end
                E: begin
                    if ((contadorCLK[7:0] == 8'b11001001))
                        reg_fstate <= S0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= E;
                end
                default: begin
                    registro <= 8'bxxxxxxxx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // tareaFSM
